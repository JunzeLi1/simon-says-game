module ssdec_ext(input logic [4:0]in, input logic enable, output logic [6:0] out);
  logic [6:0] LED [25:0];
  assign LED[5'h0] = 7'b0111111;
  assign LED[5'h1] = 7'b0000110;
  assign LED[5'h2] = 7'b1011011;
  assign LED[5'h3] = 7'b1001111;
  assign LED[5'h4] = 7'b1100110;
  assign LED[5'h5] = 7'b1101101;
  assign LED[5'h6] = 7'b1111101;
  assign LED[5'h7] = 7'b0000111;
  assign LED[5'h8] = 7'b1111111;
  assign LED[5'h9] = 7'b1100111;
  assign LED[5'ha] = 7'b1110111;
  assign LED[5'hb] = 7'b1111100;
  assign LED[5'hc] = 7'b0111001;
  assign LED[5'hd] = 7'b1011110;
  assign LED[5'he] = 7'b1111001;
  assign LED[5'hf] = 7'b1110001;
  assign LED[{1'b1, 4'h0}] = 7'b1101111;
  assign LED[{1'b1, 4'h1}] = 7'b1110110;
  assign LED[{1'b1, 4'h2}] = 7'b0010000;
  assign LED[{1'b1, 4'h3}] = 7'b0011110;
  assign LED[{1'b1, 4'h4}] = 7'b0111000;
  assign LED[{1'b1, 4'h5}] = 7'b1010100;
  assign LED[{1'b1, 4'h6}] = 7'b1010000;
  assign LED[{1'b1, 4'h7}] = 7'b1111000;
  assign LED[{1'b1, 4'h8}] = 7'b1101110;
  assign LED[{1'b1, 4'h9}] = 7'b1010011;
  assign out[6:0] = enable ? LED[in]:0;
endmodule
